// *********************************************************************
// 
// Copyright (C) 2021-20xx CrazyBird Corporation
// 
// Filename     :   bilinear_interpolation.v
// Author       :   CrazyBird
// Email        :   CrazyBirdLin@qq.com
// 
// Description  :   
// 
// Modification History
// Date         By          Version         Change Description
//----------------------------------------------------------------------
// 2021/03/27   CrazyBird   1.0             Original
// 
// *********************************************************************
module bilinear_interpolation
#(
    parameter C_SRC_IMG_WIDTH  = 12'd640    ,
    parameter C_SRC_IMG_HEIGHT = 12'd480   
    // parameter C_DST_IMG_WIDTH  = 11'd10   ,
    // parameter C_DST_IMG_HEIGHT = 11'd8    ,
    // parameter C_X_RATIO        = 16'd32768  ,           //  floor(C_SRC_IMG_WIDTH/C_DST_IMG_WIDTH*2^16)
    // parameter C_Y_RATIO        = 16'd32768              //  floor(C_SRC_IMG_HEIGHT/C_DST_IMG_HEIGHT*2^16)
)
(
    input  wire                 clk_in1         ,
    input  wire                 clk_in2         ,
    input  wire                 rst_n           ,
    
    //  Image data prepared to be processed
    input  wire                 per_img_vsync   ,       //  Prepared Image data vsync valid signal
    input  wire                 per_img_href    ,       //  Prepared Image data href vaild  signal
    input  wire     [7:0]       per_img_gray    ,       //  Prepared Image brightness input
    
    //  Image data has been processed
    output reg                  post_img_vsync  ,       //  processed Image data vsync valid signal
    output reg                  post_img_href   ,       //  processed Image data href vaild  signal
    output reg      [7:0]       post_img_gray  ,         //  processed Image brightness output

    input  wire  [11:0] c_dst_img_width,
    input  wire  [11:0] c_dst_img_height,
    output reg         [11:0]              C_DST_IMG_WIDTH,
    output reg         [11:0]              C_DST_IMG_HEIGHT
);
//----------------------------------------------------------------------

//--------------------------------my own--------------------------------------

reg                             post_img_vsync_dly;
wire                            post_img_vsync_neg;
always @(posedge clk_in2)
begin
    if(rst_n == 1'b0)
        post_img_vsync_dly <= 1'b0;
    else
        post_img_vsync_dly <= post_img_vsync;
end
assign post_img_vsync_neg = post_img_vsync_dly & ~post_img_vsync;


// c1-----

reg                             post_img_vsync_neg_c1;
always@(posedge clk_in2)
begin
    if(rst_n == 1'b0)begin
        post_img_vsync_neg_c1 =0;
    end
    else begin
        post_img_vsync_neg_c1 <=post_img_vsync_neg;
    end
end

//c1.5
reg                             post_img_vsync_neg_c1_5;
always@(posedge clk_in2)
begin
    if(rst_n == 1'b0)begin
        post_img_vsync_neg_c1_5 =0;
    end
    else begin
        post_img_vsync_neg_c1_5 <=post_img_vsync_neg_c1;
    end
end


// c2-----

reg                             post_img_vsync_neg_c2;
always@(posedge clk_in2)
begin
    if(rst_n == 1'b0)begin
        C_DST_IMG_WIDTH  <= 640;
        C_DST_IMG_HEIGHT <= 480;
    end
    else begin
        if(post_img_vsync_neg_c1_5 == 1) 
        begin
            C_DST_IMG_WIDTH  <= c_dst_img_width;
            C_DST_IMG_HEIGHT <= c_dst_img_height;
            post_img_vsync_neg_c2 <= 1;
        end
        else
        begin
            C_DST_IMG_WIDTH  <= C_DST_IMG_WIDTH;
            C_DST_IMG_HEIGHT <= C_DST_IMG_HEIGHT;
            post_img_vsync_neg_c2 <= 0;
        end
    end
end


//c3-----
reg             [26:0]          multi_tmp1_c2;
reg             [26:0]          multi_tmp2_c2;
reg                             post_img_vsync_neg_c3;

always@(posedge clk_in2)
begin
    if(rst_n == 1'b0)begin
        multi_tmp1_c2  <= 0;
        multi_tmp2_c2  <= 0;
    end
    else begin
        if(post_img_vsync_neg_c2 ==1) begin
            multi_tmp1_c2 <=(C_SRC_IMG_WIDTH <<16) ;// C_DST_IMG_WIDTH ;//  floor(C_SRC_IMG_WIDTH/C_DST_IMG_WIDTH*2^16)
            multi_tmp2_c2 <=(C_SRC_IMG_HEIGHT <<16) ;// C_DST_IMG_HEIGHT ;//  floor(C_SRC_IMG_HEIGHT/C_DST_IMG_HEIGHT*2^16)
            post_img_vsync_neg_c3 <=1;
        end
        else begin
            multi_tmp1_c2 <=multi_tmp1_c2;
            multi_tmp2_c2 <=multi_tmp2_c2;
            post_img_vsync_neg_c3 <=0;
        end
    end
end

//c4-------
reg         [18:0]              C_X_RATIO;
reg         [18:0]              C_Y_RATIO;
reg    divide_clken;
wire    rfd;
wire    rfd1;
wire   [26:0]   c_x_ratio_divide;
wire   [26:0]   c_y_ratio_divide;
always@(posedge clk_in2)
begin
    if(rst_n == 1'b0)begin
        divide_clken  <= 0; 
    end
    else begin
        if(post_img_vsync_neg_c3 ==1 && rfd ==0) begin
            divide_clken <= 1;
        end
        else if(post_img_vsync_neg_c3 ==0 && rfd ==1) begin
            divide_clken <= 0;
        end else
            divide_clken <= divide_clken;
    end
end

divider_ip ux_divider_ip(  
    .numer(multi_tmp1_c2), //  floor(C_SRC_IMG_WIDTH/C_DST_IMG_WIDTH*2^16)
    .denom(C_DST_IMG_WIDTH),
    .clken(divide_clken),
    .clk(clk_in2),
    .reset(1'b0),
    .quotient(c_x_ratio_divide),
    .remain(),
    .rfd(rfd1)

);
divider_ip uy_divider_ip(
    .numer(multi_tmp2_c2),
    .denom(C_DST_IMG_HEIGHT),
    .clken(divide_clken),
    .clk(clk_in2),
    .reset(1'b0),
    .quotient(c_y_ratio_divide),
    .remain(),
    .rfd(rfd)

);
always@(posedge clk_in2)
begin
    if(rst_n == 1'b0)begin
        C_X_RATIO  <= 65536; 
        C_Y_RATIO  <= 65536; 
    end
    else begin
        if (rfd ==1) begin
            C_X_RATIO  <= c_x_ratio_divide; 
            C_Y_RATIO  <= c_y_ratio_divide; 
        end else begin
            C_X_RATIO  <= C_X_RATIO; 
            C_Y_RATIO  <= C_Y_RATIO; 
        end
    end
end












//---------------------------end my own---------------------------------------------------



//from this ,the code is right

reg                             per_img_href_dly;

always @(posedge clk_in1)
begin
    if(rst_n == 1'b0)
        per_img_href_dly <= 1'b0;
    else
        per_img_href_dly <= per_img_href;
end

wire                            per_img_href_neg;

assign per_img_href_neg = per_img_href_dly & ~per_img_href;

reg             [10:0]          img_vs_cnt;                             //  from 0 to C_SRC_IMG_HEIGHT - 1

always @(posedge clk_in1)
begin
    if(rst_n == 1'b0)
        img_vs_cnt <= 11'b0;
    else
    begin
        if(per_img_vsync == 1'b0)
            img_vs_cnt <= 11'b0;
        else
        begin
            if(per_img_href_neg == 1'b1)
                img_vs_cnt <= img_vs_cnt + 1'b1;
            else
                img_vs_cnt <= img_vs_cnt;
        end
    end
end

reg             [10:0]          img_hs_cnt;                             //  from 0 to C_SRC_IMG_WIDTH - 1

always @(posedge clk_in1)
begin
    if(rst_n == 1'b0)
        img_hs_cnt <= 11'b0;
    else
    begin
        if((per_img_vsync == 1'b1)&&(per_img_href == 1'b1))
            img_hs_cnt <= img_hs_cnt + 1'b1;
        else
            img_hs_cnt <= 11'b0;
    end
end

//----------------------------------------------------------------------
reg             [7:0]           bram_a_wdata;

always @(posedge clk_in1)
begin
    bram_a_wdata <= per_img_gray;
end

reg             [11:0]          bram_a_waddr;

always @(posedge clk_in1)
begin
    bram_a_waddr <= {img_vs_cnt[2:1],10'b0} + img_hs_cnt;
end

reg                             bram1_a_wenb;

always @(posedge clk_in1)
begin
    if(rst_n == 1'b0)
        bram1_a_wenb <= 1'b0;
    else
        bram1_a_wenb <= per_img_vsync & per_img_href & ~img_vs_cnt[0];
end

reg                             bram2_a_wenb;

always @(posedge clk_in1)
begin
    if(rst_n == 1'b0)
        bram2_a_wenb <= 1'b0;
    else
        bram2_a_wenb <= per_img_vsync & per_img_href & img_vs_cnt[0];
end

reg             [10:0]          fifo_wdata;

always @(posedge clk_in1)
begin
    fifo_wdata <= img_vs_cnt;
end

reg                             fifo_wenb;

always @(posedge clk_in1)
begin
    if(rst_n == 1'b0)
        fifo_wenb <= 1'b0;
    else
    begin
        if((per_img_vsync == 1'b1)&&(per_img_href == 1'b1)&&(img_hs_cnt == C_SRC_IMG_WIDTH - 1'b1))
            fifo_wenb <= 1'b1;
        else
            fifo_wenb <= 1'b0;
    end
end

//----------------------------------------------------------------------
//  bram & fifo rw
reg             [11:0]          even_bram1_b_raddr;
reg             [11:0]          odd_bram1_b_raddr;
reg             [11:0]          even_bram2_b_raddr;
reg             [11:0]          odd_bram2_b_raddr;
wire            [ 7:0]          even_bram1_b_rdata;
wire            [ 7:0]          odd_bram1_b_rdata;
wire            [ 7:0]          even_bram2_b_rdata;
wire            [ 7:0]          odd_bram2_b_rdata;


// my_bram_ip    my_bram_ip_inst1 (
//     .address_a                         ( bram_a_waddr ),
//     .address_b                         ( even_bram1_b_raddr ),
//     .clock_a                           ( clk_in1 ),
//     .clock_b                           ( clk_in2 ),
//     .data_a                            ( bram_a_wdata ),
//     .data_b                            ( 8'b0 ),
//     .wren_a                            ( bram1_a_wenb ),
//     .wren_b                            ( 1'b0 ),
//     .q_a                               (  ),
//     .q_b                               ( even_bram1_b_rdata ) 
//     );

my_bram_ip  u1_my_bram_ip(
    .clk_a                             (    clk_in1                        ),
    .we_a                              (    bram1_a_wenb                   ),
    .addr_a                            (    bram_a_waddr                   ),
    .wdata_a                           (    bram_a_wdata                   ),
    .rdata_a                           (                                   ),
    .clk_b                             (    clk_in2                        ), 
    .we_b                              (    1'b0                           ),
    .addr_b                            (    even_bram1_b_raddr             ),
    .wdata_b                           (    8'b0                           ),
    .rdata_b                           (    even_bram1_b_rdata             )
);
my_bram_ip  u2_my_bram_ip(
    .clk_a                             (    clk_in1                     ),
    .we_a                              (    bram1_a_wenb                ),
    .addr_a                            (    bram_a_waddr                ),
    .wdata_a                           (    bram_a_wdata                ),
    .rdata_a                           (                                ),
    .clk_b                             (    clk_in2                     ), 
    .we_b                              (    1'b0                        ),
    .addr_b                            (    odd_bram1_b_raddr           ),
    .wdata_b                           (    8'b0                        ),
    .rdata_b                           (    odd_bram1_b_rdata           )
);
my_bram_ip  u3_my_bram_ip(
    .clk_a                             (      clk_in1                   ),
    .we_a                              (      bram2_a_wenb              ),
    .addr_a                            (      bram_a_waddr              ),
    .wdata_a                           (      bram_a_wdata              ),
    .rdata_a                           (                                ),
    .clk_b                             (      clk_in2                   ), 
    .we_b                              (      1'b0                      ),
    .addr_b                            (      even_bram2_b_raddr        ),
    .wdata_b                           (      8'b0                      ),
    .rdata_b                           (      even_bram2_b_rdata        )
);
my_bram_ip  u4_my_bram_ip(
    .clk_a                             (      clk_in1                     ),
    .we_a                              (      bram2_a_wenb                ),
    .addr_a                            (      bram_a_waddr                ),
    .wdata_a                           (      bram_a_wdata                ),
    .rdata_a                           (                                  ),
    .clk_b                             (      clk_in2                     ), 
    .we_b                              (      1'b0                        ),
    .addr_b                            (      odd_bram2_b_raddr           ),
    .wdata_b                           (      8'b0                        ),
    .rdata_b                           (      odd_bram2_b_rdata           )
);


    // my_bram_ip    my_bram_ip_inst1 (
    // .clock_a                           (   clk_in1                  ),
    // .wren_a                            (   bram1_a_wenb             ),
    // .address_a                         (   bram_a_waddr             ),
    // .data_a                            (   bram_a_wdata             ),
    // .q_a                               (                            ),
    // .clock_b                           (   clk_in2                  ),
    // .wren_b                            (   1'b0                     ),
    // .address_b                         (   even_bram1_b_raddr       ),
    // .data_b                            (   8'b0                     ),
    // .q_b                               (   even_bram1_b_rdata       ) 
    //     );
    // my_bram_ip    my_bram_ip_inst2 (
    // .clock_a                           (  clk_in1                   ),
    // .wren_a                            (  bram1_a_wenb              ),
    // .address_a                         (  bram_a_waddr              ),
    // .data_a                            (  bram_a_wdata              ),
    // .q_a                               (                            ),
    // .clock_b                           (  clk_in2                   ),
    // .wren_b                            (  1'b0                      ),
    // .address_b                         (  odd_bram1_b_raddr         ),
    // .data_b                            (  8'b0                      ),
    // .q_b                               (  odd_bram1_b_rdata         ) 
    //     );
    // my_bram_ip    my_bram_ip_inst3 (
    // .clock_a                           (   clk_in1                  ),
    // .wren_a                            (   bram2_a_wenb             ),
    // .address_a                         (   bram_a_waddr             ),
    // .data_a                            (   bram_a_wdata             ),
    // .q_a                               (                            ),
    // .clock_b                           (   clk_in2                  ),
    // .wren_b                            (   1'b0                     ),
    // .address_b                         (   even_bram2_b_raddr       ),
    // .data_b                            (   8'b0                     ),
    // .q_b                               (   even_bram2_b_rdata       ) 
    //     );
    // my_bram_ip    my_bram_ip_inst4 (
    // .clock_a                           ( clk_in1                   ),
    // .wren_a                            ( bram2_a_wenb              ),
    // .address_a                         ( bram_a_waddr              ),
    // .data_a                            ( bram_a_wdata              ),
    // .q_a                               (                           ),
    // .clock_b                           ( clk_in2                   ),
    // .wren_b                            ( 1'b0                      ),
    // .address_b                         ( odd_bram2_b_raddr         ),
    // .data_b                            ( 8'b0                      ),
    // .q_b                               ( odd_bram2_b_rdata         ) 
    //     );
    

//     my_bram_ip    my_bram_ip_inst2 (
//     .wren_a                            (bram1_a_wenb                ),
//     .wren_b                            (1'b0                        ),
//     .address_a                         (bram_a_waddr                ),
//     .data_a                            (bram_a_wdata                ),
//     .q_a                               (                            ),
//     .q_b                               (odd_bram1_b_rdata           ),
//     .address_b                         (odd_bram1_b_raddr           ),
//     .data_b                            (8'b0                        ),
//     .clock_a                           (clk_in1                     ),
//     .clock_b                           (clk_in2                     )
//         );

// my_bram_ip    my_bram_ip_inst3 (
//     .wren_a                            (bram2_a_wenb               ),
//     .wren_b                            (1'b0                       ),
//     .address_a                         (bram_a_waddr               ),
//     .data_a                            (bram_a_wdata               ),
//     .q_a                               (                           ),
//     .q_b                               (even_bram2_b_rdata         ),
//     .address_b                         (even_bram2_b_raddr         ),
//     .data_b                            (8'b0                       ),
//     .clock_a                           (clk_in1                    ),
//     .clock_b                           (clk_in2                    )
//         );


// my_bram_ip    my_bram_ip_inst4 (
//     .wren_a                            (bram2_a_wenb               ),
//     .wren_b                            (1'b0                       ),
//     .address_a                         (bram_a_waddr               ),
//     .data_a                            (bram_a_wdata               ),
//     .q_a                               (                           ),
//     .q_b                               (odd_bram2_b_rdata          ),
//     .address_b                         (odd_bram2_b_raddr          ),
//     .data_b                            (8'b0                       ),
//     .clock_a                           (clk_in1                    ),
//     .clock_b                           (clk_in2                    )
//         );
wire                            fifo_renb;
wire            [10:0]          fifo_rdata;
wire                            fifo_empty;
wire                            fifo_full;



// my_altera_fifo    my_altera_fifo_inst (
//     .aclr                              (~rst_n                    ),
//     .data                              (fifo_wdata                ),
//     .rdclk                             (clk_in2                   ),
//     .rdreq                             (fifo_renb                 ),
//     .wrclk                             (clk_in1                   ),
//     .wrreq                             (fifo_wenb                 ),
//     .q                                 (fifo_rdata                ),
//     .rdempty                           (fifo_empty                ),
//     .wrfull                            (fifo_full                 ) 
//     );

    // my_altera_fifo    my_altera_fifo_inst (
    // .aclr                              (~rst_n              ),
    // .data                              ( fifo_wdata            ),
    // .rdclk                             (  clk_in2           ),
    // .rdreq                             (   fifo_renb          ),
    // .wrclk                             (    clk_in1         ),
    // .wrreq                             (    fifo_wenb         ),
    // .q                                 (    fifo_rdata         ),
    // .rdempty                           (   fifo_empty          ),
    // .wrfull                            (    fifo_full         ) 
    // );

    asyn_fifo  u_asyn_fifo(
        .a_rst_i                           (   ~rst_n                       ), 
        .wdata                             (    fifo_wdata                  ),
        .rd_clk_i                          (     clk_in2                    ),
        .rd_en_i                           (      fifo_renb                 ),
        .wr_clk_i                          (       clk_in1                  ),
        .wr_en_i                           (       fifo_wenb                ),
        .rdata                             (       fifo_rdata               ),
        .full_o                            (      fifo_empty                ),
        .empty_o                           (       fifo_full                ),
    .almost_full_o                     (        ),
    .prog_full_o                       (        ),
    .overflow_o                        (        ),
    .wr_ack_o                          (        ),
    .almost_empty_o                    (        ),
    .underflow_o                       (        ),
    .rd_valid_o                        (        ),
    .wr_datacount_o                    (        ),
    .rst_busy                          (        ),
    .rd_datacount_o                    (        )
);


localparam S_IDLE      = 3'd0;
localparam S_Y_LOAD    = 3'd1;
localparam S_BRAM_ADDR = 3'd2;
localparam S_Y_INC     = 3'd3;
localparam S_RD_FIFO   = 3'd4;

reg             [ 2:0]          state;
reg             [26:0]          y_dec;
reg             [26:0]          x_dec;
reg             [11:0]          y_cnt;
reg             [11:0]          x_cnt;

always @(posedge clk_in2)
begin
    if(rst_n == 1'b0)
        state <= S_IDLE;
    else
    begin
        case(state)
            S_IDLE : 
            begin
                if(fifo_empty == 1'b0)
                begin
                    if((fifo_rdata != 11'b0)&&(y_cnt == C_DST_IMG_HEIGHT))
                        state <= S_RD_FIFO;
                    else
                        state <= S_Y_LOAD;
                end
                else
                    state <= S_IDLE;
            end
            S_Y_LOAD : 
            begin
                if((y_dec[26:16] + 1'b1 <= fifo_rdata)||(y_cnt == C_DST_IMG_HEIGHT - 1'b1)||((y_cnt == C_DST_IMG_HEIGHT - 2'd2)&&(C_DST_IMG_HEIGHT>=2*C_SRC_IMG_HEIGHT))||((y_cnt == C_DST_IMG_HEIGHT - 2'd3)&&(C_DST_IMG_HEIGHT>=3*C_SRC_IMG_HEIGHT))||((y_cnt == C_DST_IMG_HEIGHT - 3'd4)&&(C_DST_IMG_HEIGHT>=4*C_SRC_IMG_HEIGHT)))
                //if((y_dec[26:16] + 1'b1 <= fifo_rdata)||(y_cnt == C_DST_IMG_HEIGHT - 1'b1))
                    state <= S_BRAM_ADDR;
                else
                    state <= S_RD_FIFO;
            end
            S_BRAM_ADDR : 
            begin
                if(x_cnt == C_DST_IMG_WIDTH - 1'b1)
                    state <= S_Y_INC;
                else
                    state <= S_BRAM_ADDR;
            end
            S_Y_INC : 
            begin
                if(y_cnt == C_DST_IMG_HEIGHT - 1'b1)
                    state <= S_RD_FIFO;
                else
                    state <= S_Y_LOAD;
            end
            S_RD_FIFO : 
            begin
                state <= S_IDLE;
            end
            default : 
            begin
                state <= S_IDLE;
            end
        endcase
    end
end

assign fifo_renb = (state == S_RD_FIFO) ? 1'b1 : 1'b0;

always @(posedge clk_in2)
begin
    if(rst_n == 1'b0)
        y_dec <= 27'b0;
    else
    begin
        if((state == S_IDLE)&&(fifo_empty == 1'b0)&&(fifo_rdata == 11'b0))
            y_dec <= 27'b0;
        else if(state == S_Y_INC)
            y_dec <= y_dec + C_Y_RATIO;
        else
            y_dec <= y_dec;
    end
end

always @(posedge clk_in2)
begin
    if(rst_n == 1'b0)
        y_cnt <= 11'b0;
    else
    begin
        if((state == S_IDLE)&&(fifo_empty == 1'b0)&&(fifo_rdata == 11'b0))
            y_cnt <= 11'b0;
        else if(state == S_Y_INC)
            y_cnt <= y_cnt + 1'b1;
        else
            y_cnt <= y_cnt;
    end
end

always @(posedge clk_in2)
begin
    if(state == S_BRAM_ADDR)
        x_dec <= x_dec + C_X_RATIO;
    else
        x_dec <= 27'b0;
end

always @(posedge clk_in2)
begin
    if(state == S_BRAM_ADDR)
        x_cnt <= x_cnt + 1'b1;
    else
        x_cnt <= 11'b0;
end

//----------------------------------------------------------------------
//  c1
reg                             img_vs_c1;
reg                             debug_flag ;

always @(posedge clk_in2)
begin
    if(rst_n == 1'b0)
    begin
        img_vs_c1 <= 1'b0;
        debug_flag <= 0;
    end
    else
    begin
        if((state == S_BRAM_ADDR)&&(x_cnt == 11'b0)&&(y_cnt == 11'b0))
            img_vs_c1 <= 1'b1;
        else if((state == S_Y_INC)&&(y_cnt == C_DST_IMG_HEIGHT - 1'b1))
        begin
            img_vs_c1 <= 1'b0;
        end
        else
            img_vs_c1 <= img_vs_c1;
    end
end

reg                             img_hs_c1;

always @(posedge clk_in2)
begin
    if(rst_n == 1'b0)
        img_hs_c1 <= 1'b0;
    else
    begin
        if(state == S_BRAM_ADDR)
            img_hs_c1 <= 1'b1;
        else
            img_hs_c1 <= 1'b0;
    end
end

reg             [10:0]          x_int_c1;
reg             [10:0]          y_int_c1;
reg             [16:0]          x_fra_c1;
reg             [16:0]          inv_x_fra_c1;
reg             [16:0]          y_fra_c1;
reg             [16:0]          inv_y_fra_c1;

always @(posedge clk_in2)
begin
    x_int_c1     <= x_dec[25:16];
    y_int_c1     <= y_dec[25:16];
    x_fra_c1     <= {1'b0,x_dec[15:0]};
    inv_x_fra_c1 <= 17'h10000 - {1'b0,x_dec[15:0]};
    y_fra_c1     <= {1'b0,y_dec[15:0]};
    inv_y_fra_c1 <= 17'h10000 - {1'b0,y_dec[15:0]};
end

//----------------------------------------------------------------------
//  c2
reg                             img_vs_c2;
reg                             img_hs_c2;

always @(posedge clk_in2)
begin
    if(rst_n == 1'b0)
    begin
        img_vs_c2 <= 1'b0;
        img_hs_c2 <= 1'b0;
    end
    else
    begin
        img_vs_c2 <= img_vs_c1;
        img_hs_c2 <= img_hs_c1;
    end
end

reg             [11:0]          bram_addr_c2;
reg             [33:0]          frac_00_c2;
reg             [33:0]          frac_01_c2;
reg             [33:0]          frac_10_c2;
reg             [33:0]          frac_11_c2;
reg                             bram_mode_c2;

always @(posedge clk_in2)
begin
    bram_addr_c2 <= {y_int_c1[2:1],10'b0} + x_int_c1;
    frac_00_c2   <= inv_x_fra_c1 * inv_y_fra_c1;
    frac_01_c2   <= x_fra_c1 * inv_y_fra_c1;
    frac_10_c2   <= inv_x_fra_c1 * y_fra_c1;
    frac_11_c2   <= x_fra_c1 * y_fra_c1;
    bram_mode_c2 <= y_int_c1[0];
end

reg                             right_pixel_extand_flag_c2;
reg                             bottom_pixel_extand_flag_c2;

always @(posedge clk_in2)
begin
    if(x_int_c1 == C_SRC_IMG_WIDTH - 1'b1)
        right_pixel_extand_flag_c2 <= 1'b1;
    else
        right_pixel_extand_flag_c2 <= 1'b0;
    if(y_int_c1 == C_SRC_IMG_HEIGHT - 1'b1)
        bottom_pixel_extand_flag_c2 <= 1'b1;
    else
        bottom_pixel_extand_flag_c2 <= 1'b0;
end

//----------------------------------------------------------------------
//  c3
reg                             img_vs_c3;
reg                             img_hs_c3;

always @(posedge clk_in2)
begin
    if(rst_n == 1'b0)
    begin
        img_vs_c3 <= 1'b0;
        img_hs_c3 <= 1'b0;
    end
    else
    begin
        img_vs_c3 <= img_vs_c2;
        img_hs_c3 <= img_hs_c2;
    end
end

always @(posedge clk_in2)
begin
    if(bram_mode_c2 == 1'b0)
    begin
        even_bram1_b_raddr <= bram_addr_c2;
        odd_bram1_b_raddr  <= bram_addr_c2 + 1'b1;
        even_bram2_b_raddr <= bram_addr_c2;
        odd_bram2_b_raddr  <= bram_addr_c2 + 1'b1;
    end
    else
    begin
        even_bram1_b_raddr <= bram_addr_c2 + 11'd1024;
        odd_bram1_b_raddr  <= bram_addr_c2 + 11'd1025;
        even_bram2_b_raddr <= bram_addr_c2;
        odd_bram2_b_raddr  <= bram_addr_c2 + 1'b1;
    end
end

reg             [33:0]          frac_00_c3;
reg             [33:0]          frac_01_c3;
reg             [33:0]          frac_10_c3;
reg             [33:0]          frac_11_c3;
reg                             bram_mode_c3;
reg                             right_pixel_extand_flag_c3;
reg                             bottom_pixel_extand_flag_c3;

always @(posedge clk_in2)
begin
    frac_00_c3                  <= frac_00_c2;
    frac_01_c3                  <= frac_01_c2;
    frac_10_c3                  <= frac_10_c2;
    frac_11_c3                  <= frac_11_c2;
    bram_mode_c3                <= bram_mode_c2;
    right_pixel_extand_flag_c3  <= right_pixel_extand_flag_c2;
    bottom_pixel_extand_flag_c3 <= bottom_pixel_extand_flag_c2;
end

//----------------------------------------------------------------------
//  c4
reg                             img_vs_c4;
reg                             img_hs_c4;

always @(posedge clk_in2)
begin
    if(rst_n == 1'b0)
    begin
        img_vs_c4 <= 1'b0;
        img_hs_c4 <= 1'b0;
    end
    else
    begin
        img_vs_c4 <= img_vs_c3;
        img_hs_c4 <= img_hs_c3;
    end
end

reg             [33:0]          frac_00_c4;
reg             [33:0]          frac_01_c4;
reg             [33:0]          frac_10_c4;
reg             [33:0]          frac_11_c4;
reg                             bram_mode_c4;
reg                             right_pixel_extand_flag_c4;
reg                             bottom_pixel_extand_flag_c4;

always @(posedge clk_in2)
begin
    frac_00_c4                  <= frac_00_c3;
    frac_01_c4                  <= frac_01_c3;
    frac_10_c4                  <= frac_10_c3;
    frac_11_c4                  <= frac_11_c3;
    bram_mode_c4                <= bram_mode_c3;
    right_pixel_extand_flag_c4  <= right_pixel_extand_flag_c3;
    bottom_pixel_extand_flag_c4 <= bottom_pixel_extand_flag_c3;
end

//----------------------------------------------------------------------
//  c5
reg                             img_vs_c5;
reg                             img_hs_c5;

always @(posedge clk_in2)
begin
    if(rst_n == 1'b0)
    begin
        img_vs_c5 <= 1'b0;
        img_hs_c5 <= 1'b0;
    end
    else
    begin
        img_vs_c5 <= img_vs_c4;
        img_hs_c5 <= img_hs_c4;
    end
end

reg             [7:0]           pixel_data00_c5;
reg             [7:0]           pixel_data01_c5;
reg             [7:0]           pixel_data10_c5;
reg             [7:0]           pixel_data11_c5;

always @(posedge clk_in2)
begin
    if(bram_mode_c4 == 1'b0)
    begin
        pixel_data00_c5 <= even_bram1_b_rdata;
        pixel_data01_c5 <= odd_bram1_b_rdata;
        pixel_data10_c5 <= even_bram2_b_rdata;
        pixel_data11_c5 <= odd_bram2_b_rdata;
    end
    else
    begin
        pixel_data00_c5 <= even_bram2_b_rdata;
        pixel_data01_c5 <= odd_bram2_b_rdata;
        pixel_data10_c5 <= even_bram1_b_rdata;
        pixel_data11_c5 <= odd_bram1_b_rdata;
    end
end

reg             [33:0]          frac_00_c5;
reg             [33:0]          frac_01_c5;
reg             [33:0]          frac_10_c5;
reg             [33:0]          frac_11_c5;
reg                             right_pixel_extand_flag_c5;
reg                             bottom_pixel_extand_flag_c5;

always @(posedge clk_in2)
begin
    frac_00_c5                  <= frac_00_c4;
    frac_01_c5                  <= frac_01_c4;
    frac_10_c5                  <= frac_10_c4;
    frac_11_c5                  <= frac_11_c4;
    right_pixel_extand_flag_c5  <= right_pixel_extand_flag_c4;
    bottom_pixel_extand_flag_c5 <= bottom_pixel_extand_flag_c4;
end

//----------------------------------------------------------------------
//  c6
reg                             img_vs_c6;
reg                             img_hs_c6;

always @(posedge clk_in2)
begin
    if(rst_n == 1'b0)
    begin
        img_vs_c6 <= 1'b0;
        img_hs_c6 <= 1'b0;
    end
    else
    begin
        img_vs_c6 <= img_vs_c5;
        img_hs_c6 <= img_hs_c5;
    end
end

reg             [7:0]           pixel_data00_c6;
reg             [7:0]           pixel_data01_c6;
reg             [7:0]           pixel_data10_c6;
reg             [7:0]           pixel_data11_c6;

always @(posedge clk_in2)
begin
    case({right_pixel_extand_flag_c5,bottom_pixel_extand_flag_c5})
        2'b00 : 
        begin
            pixel_data00_c6 <= pixel_data00_c5;
            pixel_data01_c6 <= pixel_data01_c5;
            pixel_data10_c6 <= pixel_data10_c5;
            pixel_data11_c6 <= pixel_data11_c5;
        end
        2'b01 : 
        begin
            pixel_data00_c6 <= pixel_data00_c5;
            pixel_data01_c6 <= pixel_data01_c5;
            pixel_data10_c6 <= pixel_data00_c5;
            pixel_data11_c6 <= pixel_data01_c5;
        end
        2'b10 : 
        begin
            pixel_data00_c6 <= pixel_data00_c5;
            pixel_data01_c6 <= pixel_data00_c5;
            pixel_data10_c6 <= pixel_data10_c5;
            pixel_data11_c6 <= pixel_data10_c5;
        end
        2'b11 : 
        begin
            pixel_data00_c6 <= pixel_data00_c5;
            pixel_data01_c6 <= pixel_data00_c5;
            pixel_data10_c6 <= pixel_data00_c5;
            pixel_data11_c6 <= pixel_data00_c5;
        end
    endcase
end

reg             [33:0]          frac_00_c6;
reg             [33:0]          frac_01_c6;
reg             [33:0]          frac_10_c6;
reg             [33:0]          frac_11_c6;

always @(posedge clk_in2)
begin
    frac_00_c6 <= frac_00_c5;
    frac_01_c6 <= frac_01_c5;
    frac_10_c6 <= frac_10_c5;
    frac_11_c6 <= frac_11_c5;
end

//----------------------------------------------------------------------
//  c7
reg                             img_vs_c7;
reg                             img_hs_c7;

always @(posedge clk_in2)
begin
    if(rst_n == 1'b0)
    begin
        img_vs_c7 <= 1'b0;
        img_hs_c7 <= 1'b0;
    end
    else
    begin
        img_vs_c7 <= img_vs_c6;
        img_hs_c7 <= img_hs_c6;
    end
end

reg             [41:0]          gray_data00_c7;
reg             [41:0]          gray_data01_c7;
reg             [41:0]          gray_data10_c7;
reg             [41:0]          gray_data11_c7;

always @(posedge clk_in2)
begin
    gray_data00_c7 <= frac_00_c6 * pixel_data00_c6;
    gray_data01_c7 <= frac_01_c6 * pixel_data01_c6;
    gray_data10_c7 <= frac_10_c6 * pixel_data10_c6;
    gray_data11_c7 <= frac_11_c6 * pixel_data11_c6;
end

//----------------------------------------------------------------------
//  c8
reg                             img_vs_c8;
reg                             img_hs_c8;

always @(posedge clk_in2)
begin
    if(rst_n == 1'b0)
    begin
        img_vs_c8 <= 1'b0;
        img_hs_c8 <= 1'b0;
    end
    else
    begin
        img_vs_c8 <= img_vs_c7;
        img_hs_c8 <= img_hs_c7;
    end
end

reg             [42:0]          gray_data_tmp1_c8;
reg             [42:0]          gray_data_tmp2_c8;

always @(posedge clk_in2)
begin
    gray_data_tmp1_c8 <= gray_data00_c7 + gray_data01_c7;
    gray_data_tmp2_c8 <= gray_data10_c7 + gray_data11_c7;
end

//----------------------------------------------------------------------
//  c9
reg                             img_vs_c9;
reg                             img_hs_c9;

always @(posedge clk_in2)
begin
    if(rst_n == 1'b0)
    begin
        img_vs_c9 <= 1'b0;
        img_hs_c9 <= 1'b0;
    end
    else
    begin
        img_vs_c9 <= img_vs_c8;
        img_hs_c9 <= img_hs_c8;
    end
end

reg             [43:0]          gray_data_c9;

always @(posedge clk_in2)
begin
    gray_data_c9 <= gray_data_tmp1_c8 + gray_data_tmp2_c8;
end

//----------------------------------------------------------------------
//  c10
reg                             img_vs_c10;
reg                             img_hs_c10;

always @(posedge clk_in2)
begin
    if(rst_n == 1'b0)
    begin
        img_vs_c10 <= 1'b0;
        img_hs_c10 <= 1'b0;
    end
    else
    begin
        img_vs_c10 <= img_vs_c9;
        img_hs_c10 <= img_hs_c9;
    end
end

reg             [11:0]          gray_data_c10;

always @(posedge clk_in2)
begin
    gray_data_c10 <= gray_data_c9[43:32] + gray_data_c9[31];
end


//img_vs_c10�½���
reg img_vs_c10_r;
wire img_vs_c10_nagedge;
always @(posedge clk_in2)begin
    if(rst_n == 1'b0)begin
        img_vs_c10_r<=1'b0;
    end
    else begin
        img_vs_c10_r<=img_vs_c10;
    end
end

assign img_vs_c10_nagedge = img_vs_c10_r&(~img_vs_c10) ? 1'b1:1'b0;

//���ź��Ӻ�20+2������
reg [4:0] img_vs_c11_cnt;
reg img_vs_c11;
reg img_vs_c10_flag;

parameter img_vs_c11_cnt_max=5'd20;
always @(posedge clk_in2)
begin
    if(rst_n == 1'b0)
    begin
        img_vs_c11 <= 1'b0;
        img_vs_c10_flag<=1'b0;        
        img_vs_c11_cnt<=5'd0;
    end
    
    else if(img_vs_c10)begin
        img_vs_c11<=1'b1;
    end
    
    else if (img_vs_c10_nagedge)
    begin 
        img_vs_c10_flag<=1'b1;
        img_vs_c11<=1'b1;
    end
    
    else if (img_vs_c10_flag && img_vs_c11_cnt<img_vs_c11_cnt_max)
    begin
        img_vs_c11 <= 1'b1;
        img_vs_c11_cnt<=img_vs_c11_cnt+5'd1;
    end
    
    else if (img_vs_c10_flag && img_vs_c11_cnt==img_vs_c11_cnt_max)
    begin
        img_vs_c11 <= 1'b0;
        img_vs_c11_cnt<=5'd0;
        img_vs_c10_flag <= 1'b0;
    end
    
    else 
    begin
        img_vs_c11 <= 1'b0;
        img_vs_c11_cnt<=5'd0;
        img_vs_c10_flag <= 1'b0;
    end
end

//----------------------------------------------------------------------
//  signals output
always @(posedge clk_in2)
begin
    if(rst_n == 1'b0)
    begin
        post_img_vsync <= 1'b0;
        post_img_href  <= 1'b0;
    end
    else
    begin
        post_img_vsync <= (img_vs_c10||img_vs_c9||img_vs_c11);//���ź���ǰһ������//�Ӻ�20������//////////////////////////
        post_img_href  <= img_hs_c10;
    end
end

always @(posedge clk_in2)
begin
    if(gray_data_c10 > 12'd255)
        post_img_gray <= 8'd255;
    else
        post_img_gray <= gray_data_c10[7:0];
end

endmodule